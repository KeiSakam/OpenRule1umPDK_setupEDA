* Extracted by KLayout

.SUBCKT TOP VIN VOUT VDD VSS
M$1 VOUT VIN VSS VSS NCHOR1EX L=1U W=2U AS=4P AD=4P PS=8U PD=8U
M$2 VOUT VIN VDD VDD PCHOR1EX L=1U W=3.3U AS=6.6P AD=6.6P PS=10.6U PD=10.6U
.ENDS TOP
