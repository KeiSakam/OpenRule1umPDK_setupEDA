* Created by KLayout

* cell TOP
.SUBCKT TOP
* net 1 in
* net 2 out
* net 3 VDD
* net 4 VSS
* cell instance $1 r0 *1 0,0.7
X$1 3 2 1 3 Pch$1
* cell instance $2 r0 *1 -0.1,-16.6
X$2 4 2 1 4 Nch$1
.ENDS TOP

* cell Nch$1
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch$1 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,4 NMOS
M$1 2 3 1 4 NMOS L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS Nch$1

* cell Pch$1
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch$1 1 2 3 4
* device instance $1 r0 *1 2.5,6 PMOS
M$1 2 3 1 4 PMOS L=1U W=6U AS=12P AD=12P PS=16U PD=16U
.ENDS Pch$1
